`include "led_tm1637.v"
`include "led_tm1637_rom.v"
`include "spi_master.v"
